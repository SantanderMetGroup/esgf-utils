netcdf rlon_rlat {
dimensions:
	rlat = 167 ;
	rlon = 146 ;
variables:
	double lat(rlat, rlon) ;
		lat:long_name = "latitude" ;
		lat:standard_name = "latitude" ;
		lat:units = "degrees_north" ;
	double lon(rlat, rlon) ;
		lon:long_name = "longitude" ;
		lon:standard_name = "longitude" ;
		lon:units = "degrees_east" ;
	char rotated_pole ;
		rotated_pole:grid_mapping_name = "rotated_latitude_longitude" ;
		rotated_pole:grid_north_pole_latitude = 70.6 ;
		rotated_pole:grid_north_pole_longitude = -56.06 ;
	double rlon(rlon) ;
		rlon:long_name = "longitude in rotated pole grid" ;
		rlon:units = "degrees" ;
		rlon:standard_name = "grid_longitude" ;
		rlon:axis = "X" ;
	double rlat(rlat) ;
		rlat:long_name = "latitude in rotated pole grid" ;
		rlat:units = "degrees" ;
		rlat:standard_name = "grid_latitude" ;
		rlat:axis = "Y" ;

// global attributes:
		:Conventions = "CF-1.7" ;
		:title = "CORDEX South America CanESM2 Run" ;
		:contact = "meteo@unican.es" ;
		:experiment = "RCP8.5" ;
		:experiment_id = "rcp85" ;
		:driving_experiment = "CCCma-CanESM2, rcp85, r1i1p1" ;
		:driving_experiment_name = "rcp85" ;
		:driving_model_id = "CCCma-CanESM2" ;
		:driving_model_ensemble_member = "r1i1p1" ;
		:frequency = "day" ;
		:institution = "Universidad de Cantabria (Spain)" ;
		:institute_id = "UCAN" ;
		:model_id = "UCAN-WRF341I" ;
		:rcm_version_id = "v2" ;
		:project_id = "CORDEX" ;
		:CORDEX_domain = "SAM-44" ;
		:product = "output" ;
		:references = "http://www.meteo.unican.es" ;
		:ucan_run_id = "SAM044_CanESM2_altamira" ;
		:ucan_run_performance = "Altamira Supercomputer at IFCA-CSIC" ;
data:

 rlon = 143.913391113281, 144.35338973999, 144.793392181396, 
    145.233390808105, 145.673389434814, 146.113391876221, 146.55339050293, 
    146.993392944336, 147.433391571045, 147.873390197754, 148.313390731812, 
    148.753391265869, 149.193389892578, 149.633390426636, 150.073390960693, 
    150.513391494751, 150.953392028809, 151.393390655518, 151.833391189575, 
    152.273391723633, 152.713390350342, 153.153390884399, 153.593391418457, 
    154.033390045166, 154.473390579224, 154.913391113281, 155.35338973999, 
    155.793392181396, 156.233390808105, 156.673391342163, 157.113391876221, 
    157.55339050293, 157.993391036987, 158.433391571045, 158.873390197754, 
    159.313390731812, 159.753391265869, 160.193391799927, 160.633390426636, 
    161.073390960693, 161.513391494751, 161.95339012146, 162.393390655518, 
    162.833391189575, 163.273391723633, 163.713390350342, 164.153390884399, 
    164.593391418457, 165.033390045166, 165.473390579224, 165.913391113281, 
    166.353391647339, 166.793390274048, 167.233390808105, 167.673391342163, 
    168.113391876221, 168.55339050293, 168.993391036987, 169.433391571045, 
    169.873390197754, 170.313390731812, 170.753391265869, 171.193391799927, 
    171.633390426636, 172.073390960693, 172.513391494751, 172.95339012146, 
    173.393390655518, 173.833391189575, 174.273391723633, 174.713390350342, 
    175.153390884399, 175.593391418457, 176.033390045166, 176.473392486572, 
    176.913391113281, 177.35338973999, 177.793392181396, 178.233390808105, 
    178.673389434814, 179.113391876221, 179.55339050293, 179.993389129639, 
    180.433391571045, 180.873390197754, 181.31339263916, 181.753391265869, 
    182.193389892578, 182.633392333984, 183.073390960693, 183.513389587402, 
    183.953392028809, 184.393390655518, 184.833389282227, 185.273391723633, 
    185.713390350342, 186.153388977051, 186.593391418457, 187.033390045166, 
    187.473392486572, 187.913391113281, 188.35338973999, 188.793392181396, 
    189.233390808105, 189.673389434814, 190.113391876221, 190.55339050293, 
    190.993389129639, 191.433391571045, 191.873390197754, 192.31339263916, 
    192.753391265869, 193.193389892578, 193.633392333984, 194.073390960693, 
    194.513389587402, 194.953392028809, 195.393390655518, 195.833389282227, 
    196.273391723633, 196.713390350342, 197.153388977051, 197.593391418457, 
    198.033390045166, 198.473392486572, 198.913391113281, 199.35338973999, 
    199.793392181396, 200.233390808105, 200.673389434814, 201.113391876221, 
    201.55339050293, 201.993389129639, 202.433391571045, 202.873390197754, 
    203.31339263916, 203.753391265869, 204.193389892578, 204.633392333984, 
    205.073390960693, 205.513389587402, 205.953392028809, 206.393390655518, 
    206.833389282227, 207.273391723633, 207.713390350342 ;

 rlat = -38.2761535644531, -37.8361511230469, -37.3961486816406, 
    -36.9561538696289, -36.5161514282227, -36.0761489868164, 
    -35.6361541748047, -35.1961517333984, -34.7561492919922, 
    -34.3161544799805, -33.8761520385742, -33.436149597168, 
    -32.9961547851562, -32.55615234375, -32.1161499023438, -31.676155090332, 
    -31.2361526489258, -30.7961502075195, -30.3561553955078, 
    -29.9161529541016, -29.4761505126953, -29.0361518859863, 
    -28.5961532592773, -28.1561508178711, -27.7161521911621, 
    -27.2761535644531, -26.8361511230469, -26.3961524963379, 
    -25.9561538696289, -25.5161514282227, -25.0761528015137, 
    -24.6361541748047, -24.1961517333984, -23.7561531066895, 
    -23.3161506652832, -22.8761520385742, -22.4361534118652, 
    -21.996150970459, -21.55615234375, -21.116153717041, -20.6761512756348, 
    -20.2361526489258, -19.7961540222168, -19.3561515808105, 
    -18.9161529541016, -18.4761505126953, -18.0361518859863, 
    -17.5961532592773, -17.1561508178711, -16.7161521911621, 
    -16.2761535644531, -15.8361511230469, -15.3961524963379, 
    -14.9561538696289, -14.5161514282227, -14.0761528015137, 
    -13.6361541748047, -13.1961517333984, -12.7561531066895, 
    -12.3161506652832, -11.8761520385742, -11.4361534118652, 
    -10.996150970459, -10.55615234375, -10.116153717041, -9.67615127563477, 
    -9.23615264892578, -8.7961540222168, -8.35615158081055, 
    -7.91615295410156, -7.47615051269531, -7.03615188598633, 
    -6.59615325927734, -6.15615081787109, -5.71615219116211, 
    -5.27615356445312, -4.83615112304688, -4.39615249633789, 
    -3.95615386962891, -3.51615142822266, -3.07615280151367, 
    -2.63615417480469, -2.19615173339844, -1.75615310668945, 
    -1.3161506652832, -0.876152038574219, -0.436153411865234, 
    0.00384902954101562, 0.44384765625, 0.883846282958984, 1.32384872436523, 
    1.76384735107422, 2.2038459777832, 2.64384841918945, 3.08384704589844, 
    3.52384757995605, 3.96384811401367, 4.40384674072266, 4.84384727478027, 
    5.28384780883789, 5.72384834289551, 6.16384696960449, 6.60384750366211, 
    7.04384803771973, 7.48384666442871, 7.92384719848633, 8.36384773254395, 
    8.80384826660156, 9.24384689331055, 9.68384742736816, 10.1238479614258, 
    10.5638465881348, 11.0038471221924, 11.44384765625, 11.8838481903076, 
    12.3238468170166, 12.7638473510742, 13.2038478851318, 13.6438484191895, 
    14.0838470458984, 14.5238475799561, 14.9638481140137, 15.4038467407227, 
    15.8438472747803, 16.2838478088379, 16.7238483428955, 17.1638469696045, 
    17.6038475036621, 18.0438480377197, 18.4838466644287, 18.9238471984863, 
    19.3638477325439, 19.8038482666016, 20.2438468933105, 20.6838474273682, 
    21.1238479614258, 21.5638465881348, 22.0038471221924, 22.44384765625, 
    22.883846282959, 23.3238487243652, 23.7638473510742, 24.2038478851318, 
    24.6438484191895, 25.0838470458984, 25.5238475799561, 25.9638481140137, 
    26.4038467407227, 26.8438472747803, 27.2838478088379, 27.7238464355469, 
    28.1638469696045, 28.6038475036621, 29.0438480377197, 29.4838485717773, 
    29.9238471984863, 30.3638477325439, 30.8038482666016, 31.2438468933105, 
    31.6838474273682, 32.1238479614258, 32.5638465881348, 33.003849029541, 
    33.44384765625, 33.883846282959, 34.3238487243652, 34.7638473510742 ;
}
